`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 18.10.2023 19:58:00
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top(input clk_in, rst_in);
        /*
        wire ack;
        wire [31:0] data_in;
        wire [4:0] addr;
        wire cyc, stb, we;
        wire [31:0]data_out;
        wire [3:0]sel_out;
        wire sclk, miso, mosi;
        wire [31:0] ss;
        wire wb_int_out;
        */

        /*wishbone_master wishbone_master(clk_in,rst_in,ack,data_in,addr,cyc,stb,we,data_out,sel_out);
        
        spi_top spi_top(clk_in,rst_in,stb,cyc,miso,
        addr,data_out,sel_out, sclk, mosi, ack, wb_int_out, data_in, ss);
        
        spi_slave spi_slave(sclk,mosi,ss,miso);*/
endmodule
